//`timescale 1ns/10ps
`include "Single_thread.sv"
`define var_num 12'd600
`define unsat_clause_num 12'd336
`define sim_time 1000
`define dp_delay_time 1
module Single_thread_tb;
  logic clk;
  logic rst;
  logic sat;
  logic [11:0] clause_num;
  logic [10:0] mem_count_init;
  always #5 clk = ~clk;
  integer fout,funsat;
 
  Single_thread s(
    .clk(clk),
    .rst(rst),
	.boot(1'b0),
	.clause_num(clause_num),
	.mem_count_init(mem_count_init),
    .sat(sat)
  );
  
  
  
  initial begin
    clk = 1'b0;
    rst = 1'b1;
	clause_num = `var_num;
	mem_count_init = 12'd336//`unsat_clause_num;
    #10
	rst = 1'b0;
	s.tt.AT.address_mem[0] = 11'bz;
    $readmemh("../addr.dat",s.tt.AT.address_mem,1);
	$readmemb("../mask.dat",s.tt.AT.Mask_mem,1);
	$readmemh("../clause_table.dat",s.tt.CT.mem,0);
	$readmemb("../true_value.dat",s.tt.cr.eva2.var_table,0);
	$readmemb("../true_value.dat",s.pe.evaluator2.var_table,0);
   // $readmemb("../true_value.dat",s.pe.idle_check.var_table,0);	
	$readmemh("../unsatisfied_clause.dat",s.pe.ucb.mem,0);
    
  end

  initial begin
    $fsdbDumpfile("Single_thread.fsdb");
    $fsdbDumpvars(0,Single_thread_tb);
	
	fout = $fopen("value.out","w");
	funsat = $fopen("unsat.out","w");
	/*for(int i=0;i<3000;++i) begin
	  #10 
	    if(sat & s.tt.cr.sat == 1'b1) begin
		  print_result();
		  $finish;
		end
	end
	*/
  end
  
  initial begin
    #`sim_time
	print_result();
    $finish;
  end
  
  initial begin
    s.tt.cr.share_memory= 600'b0;
    s.tt.cr.assign_memory= 600'b0;
    #`dp_delay_time
s.tt.cr.share_memory[1]= 1'b0;
s.tt.cr.assign_memory[1]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[2]= 1'b1;
s.tt.cr.assign_memory[2]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[3]= 1'b0;
s.tt.cr.assign_memory[3]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[4]= 1'b1;
s.tt.cr.assign_memory[4]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[5]= 1'b0;
s.tt.cr.assign_memory[5]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[6]= 1'b0;
s.tt.cr.assign_memory[6]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[7]= 1'b1;
s.tt.cr.assign_memory[7]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[8]= 1'b0;
s.tt.cr.assign_memory[8]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[9]= 1'b1;
s.tt.cr.assign_memory[9]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[10]= 1'b1;
s.tt.cr.assign_memory[10]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[11]= 1'b1;
s.tt.cr.assign_memory[11]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[12]= 1'b1;
s.tt.cr.assign_memory[12]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[13]= 1'b1;
s.tt.cr.assign_memory[13]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[14]= 1'b0;
s.tt.cr.assign_memory[14]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[15]= 1'b1;
s.tt.cr.assign_memory[15]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[16]= 1'b1;
s.tt.cr.assign_memory[16]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[17]= 1'b1;
s.tt.cr.assign_memory[17]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[18]= 1'b1;
s.tt.cr.assign_memory[18]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[19]= 1'b1;
s.tt.cr.assign_memory[19]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[20]= 1'b0;
s.tt.cr.assign_memory[20]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[21]= 1'b0;
s.tt.cr.assign_memory[21]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[22]= 1'b0;
s.tt.cr.assign_memory[22]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[23]= 1'b1;
s.tt.cr.assign_memory[23]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[24]= 1'b1;
s.tt.cr.assign_memory[24]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[25]= 1'b1;
s.tt.cr.assign_memory[25]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[26]= 1'b0;
s.tt.cr.assign_memory[26]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[27]= 1'b0;
s.tt.cr.assign_memory[27]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[28]= 1'b1;
s.tt.cr.assign_memory[28]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[29]= 1'b0;
s.tt.cr.assign_memory[29]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[30]= 1'b0;
s.tt.cr.assign_memory[30]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[31]= 1'b1;
s.tt.cr.assign_memory[31]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[32]= 1'b0;
s.tt.cr.assign_memory[32]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[33]= 1'b1;
s.tt.cr.assign_memory[33]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[34]= 1'b1;
s.tt.cr.assign_memory[34]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[35]= 1'b1;
s.tt.cr.assign_memory[35]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[36]= 1'b1;
s.tt.cr.assign_memory[36]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[37]= 1'b0;
s.tt.cr.assign_memory[37]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[38]= 1'b1;
s.tt.cr.assign_memory[38]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[39]= 1'b1;
s.tt.cr.assign_memory[39]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[40]= 1'b0;
s.tt.cr.assign_memory[40]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[41]= 1'b1;
s.tt.cr.assign_memory[41]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[42]= 1'b0;
s.tt.cr.assign_memory[42]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[43]= 1'b1;
s.tt.cr.assign_memory[43]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[44]= 1'b0;
s.tt.cr.assign_memory[44]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[45]= 1'b1;
s.tt.cr.assign_memory[45]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[46]= 1'b0;
s.tt.cr.assign_memory[46]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[47]= 1'b1;
s.tt.cr.assign_memory[47]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[48]= 1'b1;
s.tt.cr.assign_memory[48]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[49]= 1'b0;
s.tt.cr.assign_memory[49]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[50]= 1'b0;
s.tt.cr.assign_memory[50]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[51]= 1'b1;
s.tt.cr.assign_memory[51]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[52]= 1'b0;
s.tt.cr.assign_memory[52]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[53]= 1'b0;
s.tt.cr.assign_memory[53]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[54]= 1'b1;
s.tt.cr.assign_memory[54]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[55]= 1'b0;
s.tt.cr.assign_memory[55]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[56]= 1'b1;
s.tt.cr.assign_memory[56]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[57]= 1'b1;
s.tt.cr.assign_memory[57]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[58]= 1'b1;
s.tt.cr.assign_memory[58]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[59]= 1'b1;
s.tt.cr.assign_memory[59]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[60]= 1'b0;
s.tt.cr.assign_memory[60]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[61]= 1'b1;
s.tt.cr.assign_memory[61]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[62]= 1'b0;
s.tt.cr.assign_memory[62]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[63]= 1'b0;
s.tt.cr.assign_memory[63]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[64]= 1'b1;
s.tt.cr.assign_memory[64]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[65]= 1'b1;
s.tt.cr.assign_memory[65]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[66]= 1'b0;
s.tt.cr.assign_memory[66]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[67]= 1'b1;
s.tt.cr.assign_memory[67]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[68]= 1'b1;
s.tt.cr.assign_memory[68]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[69]= 1'b0;
s.tt.cr.assign_memory[69]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[70]= 1'b0;
s.tt.cr.assign_memory[70]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[71]= 1'b0;
s.tt.cr.assign_memory[71]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[72]= 1'b0;
s.tt.cr.assign_memory[72]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[73]= 1'b1;
s.tt.cr.assign_memory[73]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[74]= 1'b0;
s.tt.cr.assign_memory[74]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[75]= 1'b1;
s.tt.cr.assign_memory[75]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[76]= 1'b0;
s.tt.cr.assign_memory[76]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[77]= 1'b0;
s.tt.cr.assign_memory[77]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[78]= 1'b1;
s.tt.cr.assign_memory[78]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[79]= 1'b1;
s.tt.cr.assign_memory[79]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[80]= 1'b1;
s.tt.cr.assign_memory[80]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[81]= 1'b0;
s.tt.cr.assign_memory[81]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[82]= 1'b1;
s.tt.cr.assign_memory[82]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[83]= 1'b0;
s.tt.cr.assign_memory[83]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[84]= 1'b1;
s.tt.cr.assign_memory[84]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[85]= 1'b1;
s.tt.cr.assign_memory[85]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[86]= 1'b1;
s.tt.cr.assign_memory[86]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[87]= 1'b0;
s.tt.cr.assign_memory[87]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[88]= 1'b1;
s.tt.cr.assign_memory[88]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[89]= 1'b1;
s.tt.cr.assign_memory[89]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[90]= 1'b0;
s.tt.cr.assign_memory[90]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[91]= 1'b0;
s.tt.cr.assign_memory[91]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[92]= 1'b0;
s.tt.cr.assign_memory[92]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[93]= 1'b1;
s.tt.cr.assign_memory[93]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[94]= 1'b1;
s.tt.cr.assign_memory[94]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[95]= 1'b0;
s.tt.cr.assign_memory[95]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[96]= 1'b1;
s.tt.cr.assign_memory[96]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[97]= 1'b1;
s.tt.cr.assign_memory[97]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[98]= 1'b0;
s.tt.cr.assign_memory[98]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[99]= 1'b1;
s.tt.cr.assign_memory[99]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[100]= 1'b0;
s.tt.cr.assign_memory[100]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[101]= 1'b1;
s.tt.cr.assign_memory[101]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[102]= 1'b1;
s.tt.cr.assign_memory[102]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[103]= 1'b1;
s.tt.cr.assign_memory[103]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[104]= 1'b0;
s.tt.cr.assign_memory[104]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[105]= 1'b0;
s.tt.cr.assign_memory[105]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[106]= 1'b1;
s.tt.cr.assign_memory[106]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[107]= 1'b1;
s.tt.cr.assign_memory[107]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[108]= 1'b1;
s.tt.cr.assign_memory[108]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[109]= 1'b0;
s.tt.cr.assign_memory[109]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[110]= 1'b1;
s.tt.cr.assign_memory[110]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[111]= 1'b0;
s.tt.cr.assign_memory[111]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[112]= 1'b0;
s.tt.cr.assign_memory[112]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[113]= 1'b1;
s.tt.cr.assign_memory[113]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[114]= 1'b0;
s.tt.cr.assign_memory[114]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[115]= 1'b1;
s.tt.cr.assign_memory[115]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[116]= 1'b1;
s.tt.cr.assign_memory[116]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[117]= 1'b1;
s.tt.cr.assign_memory[117]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[118]= 1'b0;
s.tt.cr.assign_memory[118]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[119]= 1'b0;
s.tt.cr.assign_memory[119]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[120]= 1'b0;
s.tt.cr.assign_memory[120]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[121]= 1'b1;
s.tt.cr.assign_memory[121]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[122]= 1'b1;
s.tt.cr.assign_memory[122]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[123]= 1'b0;
s.tt.cr.assign_memory[123]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[124]= 1'b1;
s.tt.cr.assign_memory[124]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[125]= 1'b0;
s.tt.cr.assign_memory[125]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[126]= 1'b0;
s.tt.cr.assign_memory[126]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[127]= 1'b1;
s.tt.cr.assign_memory[127]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[128]= 1'b0;
s.tt.cr.assign_memory[128]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[129]= 1'b0;
s.tt.cr.assign_memory[129]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[130]= 1'b0;
s.tt.cr.assign_memory[130]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[131]= 1'b0;
s.tt.cr.assign_memory[131]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[132]= 1'b1;
s.tt.cr.assign_memory[132]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[133]= 1'b1;
s.tt.cr.assign_memory[133]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[134]= 1'b0;
s.tt.cr.assign_memory[134]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[135]= 1'b1;
s.tt.cr.assign_memory[135]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[136]= 1'b1;
s.tt.cr.assign_memory[136]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[137]= 1'b0;
s.tt.cr.assign_memory[137]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[138]= 1'b1;
s.tt.cr.assign_memory[138]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[139]= 1'b0;
s.tt.cr.assign_memory[139]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[140]= 1'b0;
s.tt.cr.assign_memory[140]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[141]= 1'b1;
s.tt.cr.assign_memory[141]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[142]= 1'b1;
s.tt.cr.assign_memory[142]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[143]= 1'b0;
s.tt.cr.assign_memory[143]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[144]= 1'b1;
s.tt.cr.assign_memory[144]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[145]= 1'b1;
s.tt.cr.assign_memory[145]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[146]= 1'b0;
s.tt.cr.assign_memory[146]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[147]= 1'b1;
s.tt.cr.assign_memory[147]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[148]= 1'b0;
s.tt.cr.assign_memory[148]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[149]= 1'b0;
s.tt.cr.assign_memory[149]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[150]= 1'b1;
s.tt.cr.assign_memory[150]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[151]= 1'b1;
s.tt.cr.assign_memory[151]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[152]= 1'b0;
s.tt.cr.assign_memory[152]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[153]= 1'b1;
s.tt.cr.assign_memory[153]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[154]= 1'b1;
s.tt.cr.assign_memory[154]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[155]= 1'b0;
s.tt.cr.assign_memory[155]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[156]= 1'b0;
s.tt.cr.assign_memory[156]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[157]= 1'b1;
s.tt.cr.assign_memory[157]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[158]= 1'b0;
s.tt.cr.assign_memory[158]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[159]= 1'b1;
s.tt.cr.assign_memory[159]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[160]= 1'b0;
s.tt.cr.assign_memory[160]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[161]= 1'b1;
s.tt.cr.assign_memory[161]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[162]= 1'b0;
s.tt.cr.assign_memory[162]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[163]= 1'b0;
s.tt.cr.assign_memory[163]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[164]= 1'b1;
s.tt.cr.assign_memory[164]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[165]= 1'b1;
s.tt.cr.assign_memory[165]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[166]= 1'b1;
s.tt.cr.assign_memory[166]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[167]= 1'b1;
s.tt.cr.assign_memory[167]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[168]= 1'b1;
s.tt.cr.assign_memory[168]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[169]= 1'b1;
s.tt.cr.assign_memory[169]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[170]= 1'b0;
s.tt.cr.assign_memory[170]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[171]= 1'b0;
s.tt.cr.assign_memory[171]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[172]= 1'b1;
s.tt.cr.assign_memory[172]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[173]= 1'b0;
s.tt.cr.assign_memory[173]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[174]= 1'b0;
s.tt.cr.assign_memory[174]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[175]= 1'b1;
s.tt.cr.assign_memory[175]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[176]= 1'b1;
s.tt.cr.assign_memory[176]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[177]= 1'b1;
s.tt.cr.assign_memory[177]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[178]= 1'b1;
s.tt.cr.assign_memory[178]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[179]= 1'b1;
s.tt.cr.assign_memory[179]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[180]= 1'b1;
s.tt.cr.assign_memory[180]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[181]= 1'b0;
s.tt.cr.assign_memory[181]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[182]= 1'b1;
s.tt.cr.assign_memory[182]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[183]= 1'b1;
s.tt.cr.assign_memory[183]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[184]= 1'b0;
s.tt.cr.assign_memory[184]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[185]= 1'b1;
s.tt.cr.assign_memory[185]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[186]= 1'b1;
s.tt.cr.assign_memory[186]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[187]= 1'b0;
s.tt.cr.assign_memory[187]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[188]= 1'b0;
s.tt.cr.assign_memory[188]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[189]= 1'b1;
s.tt.cr.assign_memory[189]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[190]= 1'b0;
s.tt.cr.assign_memory[190]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[191]= 1'b0;
s.tt.cr.assign_memory[191]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[192]= 1'b0;
s.tt.cr.assign_memory[192]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[193]= 1'b0;
s.tt.cr.assign_memory[193]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[194]= 1'b1;
s.tt.cr.assign_memory[194]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[195]= 1'b1;
s.tt.cr.assign_memory[195]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[196]= 1'b0;
s.tt.cr.assign_memory[196]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[197]= 1'b0;
s.tt.cr.assign_memory[197]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[198]= 1'b1;
s.tt.cr.assign_memory[198]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[199]= 1'b0;
s.tt.cr.assign_memory[199]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[200]= 1'b0;
s.tt.cr.assign_memory[200]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[201]= 1'b1;
s.tt.cr.assign_memory[201]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[202]= 1'b0;
s.tt.cr.assign_memory[202]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[203]= 1'b1;
s.tt.cr.assign_memory[203]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[204]= 1'b1;
s.tt.cr.assign_memory[204]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[205]= 1'b0;
s.tt.cr.assign_memory[205]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[206]= 1'b1;
s.tt.cr.assign_memory[206]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[207]= 1'b0;
s.tt.cr.assign_memory[207]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[208]= 1'b0;
s.tt.cr.assign_memory[208]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[209]= 1'b1;
s.tt.cr.assign_memory[209]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[210]= 1'b0;
s.tt.cr.assign_memory[210]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[211]= 1'b0;
s.tt.cr.assign_memory[211]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[212]= 1'b1;
s.tt.cr.assign_memory[212]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[213]= 1'b1;
s.tt.cr.assign_memory[213]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[214]= 1'b0;
s.tt.cr.assign_memory[214]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[215]= 1'b1;
s.tt.cr.assign_memory[215]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[216]= 1'b0;
s.tt.cr.assign_memory[216]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[217]= 1'b0;
s.tt.cr.assign_memory[217]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[218]= 1'b1;
s.tt.cr.assign_memory[218]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[219]= 1'b1;
s.tt.cr.assign_memory[219]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[220]= 1'b0;
s.tt.cr.assign_memory[220]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[221]= 1'b0;
s.tt.cr.assign_memory[221]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[222]= 1'b0;
s.tt.cr.assign_memory[222]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[223]= 1'b0;
s.tt.cr.assign_memory[223]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[224]= 1'b0;
s.tt.cr.assign_memory[224]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[225]= 1'b0;
s.tt.cr.assign_memory[225]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[226]= 1'b1;
s.tt.cr.assign_memory[226]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[227]= 1'b0;
s.tt.cr.assign_memory[227]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[228]= 1'b0;
s.tt.cr.assign_memory[228]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[229]= 1'b1;
s.tt.cr.assign_memory[229]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[230]= 1'b0;
s.tt.cr.assign_memory[230]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[231]= 1'b1;
s.tt.cr.assign_memory[231]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[232]= 1'b1;
s.tt.cr.assign_memory[232]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[233]= 1'b0;
s.tt.cr.assign_memory[233]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[234]= 1'b1;
s.tt.cr.assign_memory[234]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[235]= 1'b0;
s.tt.cr.assign_memory[235]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[236]= 1'b0;
s.tt.cr.assign_memory[236]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[237]= 1'b0;
s.tt.cr.assign_memory[237]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[238]= 1'b1;
s.tt.cr.assign_memory[238]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[239]= 1'b0;
s.tt.cr.assign_memory[239]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[240]= 1'b0;
s.tt.cr.assign_memory[240]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[241]= 1'b0;
s.tt.cr.assign_memory[241]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[242]= 1'b0;
s.tt.cr.assign_memory[242]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[243]= 1'b0;
s.tt.cr.assign_memory[243]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[244]= 1'b1;
s.tt.cr.assign_memory[244]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[245]= 1'b0;
s.tt.cr.assign_memory[245]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[246]= 1'b0;
s.tt.cr.assign_memory[246]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[247]= 1'b1;
s.tt.cr.assign_memory[247]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[248]= 1'b0;
s.tt.cr.assign_memory[248]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[249]= 1'b0;
s.tt.cr.assign_memory[249]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[250]= 1'b1;
s.tt.cr.assign_memory[250]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[251]= 1'b0;
s.tt.cr.assign_memory[251]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[252]= 1'b1;
s.tt.cr.assign_memory[252]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[253]= 1'b0;
s.tt.cr.assign_memory[253]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[254]= 1'b0;
s.tt.cr.assign_memory[254]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[255]= 1'b0;
s.tt.cr.assign_memory[255]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[256]= 1'b0;
s.tt.cr.assign_memory[256]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[257]= 1'b0;
s.tt.cr.assign_memory[257]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[258]= 1'b0;
s.tt.cr.assign_memory[258]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[259]= 1'b1;
s.tt.cr.assign_memory[259]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[260]= 1'b0;
s.tt.cr.assign_memory[260]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[261]= 1'b0;
s.tt.cr.assign_memory[261]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[262]= 1'b0;
s.tt.cr.assign_memory[262]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[263]= 1'b0;
s.tt.cr.assign_memory[263]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[264]= 1'b1;
s.tt.cr.assign_memory[264]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[265]= 1'b1;
s.tt.cr.assign_memory[265]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[266]= 1'b0;
s.tt.cr.assign_memory[266]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[267]= 1'b1;
s.tt.cr.assign_memory[267]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[268]= 1'b0;
s.tt.cr.assign_memory[268]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[269]= 1'b1;
s.tt.cr.assign_memory[269]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[270]= 1'b1;
s.tt.cr.assign_memory[270]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[271]= 1'b1;
s.tt.cr.assign_memory[271]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[272]= 1'b1;
s.tt.cr.assign_memory[272]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[273]= 1'b0;
s.tt.cr.assign_memory[273]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[274]= 1'b1;
s.tt.cr.assign_memory[274]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[275]= 1'b0;
s.tt.cr.assign_memory[275]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[276]= 1'b0;
s.tt.cr.assign_memory[276]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[277]= 1'b0;
s.tt.cr.assign_memory[277]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[278]= 1'b0;
s.tt.cr.assign_memory[278]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[279]= 1'b0;
s.tt.cr.assign_memory[279]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[280]= 1'b1;
s.tt.cr.assign_memory[280]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[281]= 1'b0;
s.tt.cr.assign_memory[281]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[282]= 1'b1;
s.tt.cr.assign_memory[282]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[283]= 1'b0;
s.tt.cr.assign_memory[283]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[284]= 1'b0;
s.tt.cr.assign_memory[284]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[285]= 1'b1;
s.tt.cr.assign_memory[285]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[286]= 1'b0;
s.tt.cr.assign_memory[286]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[287]= 1'b1;
s.tt.cr.assign_memory[287]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[288]= 1'b0;
s.tt.cr.assign_memory[288]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[289]= 1'b0;
s.tt.cr.assign_memory[289]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[290]= 1'b1;
s.tt.cr.assign_memory[290]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[291]= 1'b0;
s.tt.cr.assign_memory[291]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[292]= 1'b1;
s.tt.cr.assign_memory[292]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[293]= 1'b1;
s.tt.cr.assign_memory[293]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[294]= 1'b0;
s.tt.cr.assign_memory[294]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[295]= 1'b0;
s.tt.cr.assign_memory[295]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[296]= 1'b0;
s.tt.cr.assign_memory[296]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[297]= 1'b0;
s.tt.cr.assign_memory[297]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[298]= 1'b0;
s.tt.cr.assign_memory[298]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[299]= 1'b0;
s.tt.cr.assign_memory[299]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[300]= 1'b0;
s.tt.cr.assign_memory[300]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[301]= 1'b1;
s.tt.cr.assign_memory[301]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[302]= 1'b1;
s.tt.cr.assign_memory[302]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[303]= 1'b0;
s.tt.cr.assign_memory[303]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[304]= 1'b1;
s.tt.cr.assign_memory[304]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[305]= 1'b0;
s.tt.cr.assign_memory[305]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[306]= 1'b1;
s.tt.cr.assign_memory[306]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[307]= 1'b0;
s.tt.cr.assign_memory[307]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[308]= 1'b0;
s.tt.cr.assign_memory[308]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[309]= 1'b1;
s.tt.cr.assign_memory[309]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[310]= 1'b0;
s.tt.cr.assign_memory[310]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[311]= 1'b0;
s.tt.cr.assign_memory[311]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[312]= 1'b0;
s.tt.cr.assign_memory[312]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[313]= 1'b0;
s.tt.cr.assign_memory[313]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[314]= 1'b0;
s.tt.cr.assign_memory[314]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[315]= 1'b0;
s.tt.cr.assign_memory[315]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[316]= 1'b1;
s.tt.cr.assign_memory[316]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[317]= 1'b1;
s.tt.cr.assign_memory[317]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[318]= 1'b0;
s.tt.cr.assign_memory[318]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[319]= 1'b1;
s.tt.cr.assign_memory[319]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[320]= 1'b1;
s.tt.cr.assign_memory[320]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[321]= 1'b1;
s.tt.cr.assign_memory[321]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[322]= 1'b1;
s.tt.cr.assign_memory[322]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[323]= 1'b0;
s.tt.cr.assign_memory[323]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[324]= 1'b1;
s.tt.cr.assign_memory[324]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[325]= 1'b0;
s.tt.cr.assign_memory[325]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[326]= 1'b0;
s.tt.cr.assign_memory[326]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[327]= 1'b0;
s.tt.cr.assign_memory[327]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[328]= 1'b0;
s.tt.cr.assign_memory[328]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[329]= 1'b0;
s.tt.cr.assign_memory[329]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[330]= 1'b0;
s.tt.cr.assign_memory[330]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[331]= 1'b1;
s.tt.cr.assign_memory[331]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[332]= 1'b1;
s.tt.cr.assign_memory[332]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[333]= 1'b1;
s.tt.cr.assign_memory[333]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[334]= 1'b1;
s.tt.cr.assign_memory[334]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[335]= 1'b1;
s.tt.cr.assign_memory[335]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[336]= 1'b0;
s.tt.cr.assign_memory[336]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[337]= 1'b0;
s.tt.cr.assign_memory[337]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[338]= 1'b1;
s.tt.cr.assign_memory[338]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[339]= 1'b0;
s.tt.cr.assign_memory[339]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[340]= 1'b0;
s.tt.cr.assign_memory[340]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[341]= 1'b1;
s.tt.cr.assign_memory[341]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[342]= 1'b1;
s.tt.cr.assign_memory[342]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[343]= 1'b1;
s.tt.cr.assign_memory[343]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[344]= 1'b1;
s.tt.cr.assign_memory[344]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[345]= 1'b0;
s.tt.cr.assign_memory[345]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[346]= 1'b0;
s.tt.cr.assign_memory[346]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[347]= 1'b1;
s.tt.cr.assign_memory[347]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[348]= 1'b0;
s.tt.cr.assign_memory[348]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[349]= 1'b0;
s.tt.cr.assign_memory[349]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[350]= 1'b1;
s.tt.cr.assign_memory[350]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[351]= 1'b0;
s.tt.cr.assign_memory[351]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[352]= 1'b0;
s.tt.cr.assign_memory[352]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[353]= 1'b0;
s.tt.cr.assign_memory[353]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[354]= 1'b0;
s.tt.cr.assign_memory[354]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[355]= 1'b1;
s.tt.cr.assign_memory[355]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[356]= 1'b1;
s.tt.cr.assign_memory[356]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[357]= 1'b1;
s.tt.cr.assign_memory[357]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[358]= 1'b0;
s.tt.cr.assign_memory[358]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[359]= 1'b1;
s.tt.cr.assign_memory[359]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[360]= 1'b1;
s.tt.cr.assign_memory[360]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[361]= 1'b0;
s.tt.cr.assign_memory[361]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[362]= 1'b1;
s.tt.cr.assign_memory[362]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[363]= 1'b1;
s.tt.cr.assign_memory[363]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[364]= 1'b0;
s.tt.cr.assign_memory[364]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[365]= 1'b0;
s.tt.cr.assign_memory[365]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[366]= 1'b1;
s.tt.cr.assign_memory[366]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[367]= 1'b1;
s.tt.cr.assign_memory[367]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[368]= 1'b0;
s.tt.cr.assign_memory[368]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[369]= 1'b0;
s.tt.cr.assign_memory[369]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[370]= 1'b1;
s.tt.cr.assign_memory[370]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[371]= 1'b0;
s.tt.cr.assign_memory[371]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[372]= 1'b0;
s.tt.cr.assign_memory[372]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[373]= 1'b0;
s.tt.cr.assign_memory[373]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[374]= 1'b0;
s.tt.cr.assign_memory[374]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[375]= 1'b1;
s.tt.cr.assign_memory[375]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[376]= 1'b1;
s.tt.cr.assign_memory[376]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[377]= 1'b1;
s.tt.cr.assign_memory[377]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[378]= 1'b1;
s.tt.cr.assign_memory[378]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[379]= 1'b0;
s.tt.cr.assign_memory[379]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[380]= 1'b0;
s.tt.cr.assign_memory[380]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[381]= 1'b1;
s.tt.cr.assign_memory[381]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[382]= 1'b1;
s.tt.cr.assign_memory[382]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[383]= 1'b0;
s.tt.cr.assign_memory[383]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[384]= 1'b0;
s.tt.cr.assign_memory[384]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[385]= 1'b0;
s.tt.cr.assign_memory[385]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[386]= 1'b0;
s.tt.cr.assign_memory[386]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[387]= 1'b1;
s.tt.cr.assign_memory[387]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[388]= 1'b1;
s.tt.cr.assign_memory[388]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[389]= 1'b0;
s.tt.cr.assign_memory[389]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[390]= 1'b1;
s.tt.cr.assign_memory[390]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[391]= 1'b0;
s.tt.cr.assign_memory[391]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[392]= 1'b1;
s.tt.cr.assign_memory[392]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[393]= 1'b0;
s.tt.cr.assign_memory[393]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[394]= 1'b1;
s.tt.cr.assign_memory[394]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[395]= 1'b1;
s.tt.cr.assign_memory[395]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[396]= 1'b1;
s.tt.cr.assign_memory[396]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[397]= 1'b1;
s.tt.cr.assign_memory[397]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[398]= 1'b0;
s.tt.cr.assign_memory[398]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[399]= 1'b1;
s.tt.cr.assign_memory[399]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[400]= 1'b0;
s.tt.cr.assign_memory[400]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[401]= 1'b0;
s.tt.cr.assign_memory[401]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[402]= 1'b1;
s.tt.cr.assign_memory[402]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[403]= 1'b1;
s.tt.cr.assign_memory[403]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[404]= 1'b1;
s.tt.cr.assign_memory[404]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[405]= 1'b1;
s.tt.cr.assign_memory[405]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[406]= 1'b1;
s.tt.cr.assign_memory[406]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[407]= 1'b1;
s.tt.cr.assign_memory[407]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[408]= 1'b0;
s.tt.cr.assign_memory[408]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[409]= 1'b1;
s.tt.cr.assign_memory[409]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[410]= 1'b0;
s.tt.cr.assign_memory[410]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[411]= 1'b1;
s.tt.cr.assign_memory[411]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[412]= 1'b0;
s.tt.cr.assign_memory[412]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[413]= 1'b0;
s.tt.cr.assign_memory[413]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[414]= 1'b0;
s.tt.cr.assign_memory[414]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[415]= 1'b0;
s.tt.cr.assign_memory[415]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[416]= 1'b1;
s.tt.cr.assign_memory[416]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[417]= 1'b1;
s.tt.cr.assign_memory[417]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[418]= 1'b0;
s.tt.cr.assign_memory[418]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[419]= 1'b0;
s.tt.cr.assign_memory[419]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[420]= 1'b0;
s.tt.cr.assign_memory[420]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[421]= 1'b1;
s.tt.cr.assign_memory[421]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[422]= 1'b0;
s.tt.cr.assign_memory[422]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[423]= 1'b0;
s.tt.cr.assign_memory[423]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[424]= 1'b0;
s.tt.cr.assign_memory[424]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[425]= 1'b0;
s.tt.cr.assign_memory[425]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[426]= 1'b1;
s.tt.cr.assign_memory[426]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[427]= 1'b0;
s.tt.cr.assign_memory[427]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[428]= 1'b0;
s.tt.cr.assign_memory[428]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[429]= 1'b0;
s.tt.cr.assign_memory[429]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[430]= 1'b1;
s.tt.cr.assign_memory[430]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[431]= 1'b1;
s.tt.cr.assign_memory[431]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[432]= 1'b1;
s.tt.cr.assign_memory[432]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[433]= 1'b1;
s.tt.cr.assign_memory[433]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[434]= 1'b0;
s.tt.cr.assign_memory[434]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[435]= 1'b1;
s.tt.cr.assign_memory[435]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[436]= 1'b0;
s.tt.cr.assign_memory[436]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[437]= 1'b1;
s.tt.cr.assign_memory[437]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[438]= 1'b1;
s.tt.cr.assign_memory[438]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[439]= 1'b1;
s.tt.cr.assign_memory[439]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[440]= 1'b0;
s.tt.cr.assign_memory[440]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[441]= 1'b0;
s.tt.cr.assign_memory[441]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[442]= 1'b1;
s.tt.cr.assign_memory[442]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[443]= 1'b1;
s.tt.cr.assign_memory[443]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[444]= 1'b0;
s.tt.cr.assign_memory[444]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[445]= 1'b0;
s.tt.cr.assign_memory[445]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[446]= 1'b1;
s.tt.cr.assign_memory[446]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[447]= 1'b0;
s.tt.cr.assign_memory[447]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[448]= 1'b1;
s.tt.cr.assign_memory[448]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[449]= 1'b0;
s.tt.cr.assign_memory[449]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[450]= 1'b1;
s.tt.cr.assign_memory[450]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[451]= 1'b0;
s.tt.cr.assign_memory[451]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[452]= 1'b0;
s.tt.cr.assign_memory[452]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[453]= 1'b0;
s.tt.cr.assign_memory[453]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[454]= 1'b1;
s.tt.cr.assign_memory[454]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[455]= 1'b0;
s.tt.cr.assign_memory[455]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[456]= 1'b0;
s.tt.cr.assign_memory[456]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[457]= 1'b1;
s.tt.cr.assign_memory[457]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[458]= 1'b0;
s.tt.cr.assign_memory[458]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[459]= 1'b1;
s.tt.cr.assign_memory[459]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[460]= 1'b0;
s.tt.cr.assign_memory[460]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[461]= 1'b1;
s.tt.cr.assign_memory[461]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[462]= 1'b0;
s.tt.cr.assign_memory[462]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[463]= 1'b1;
s.tt.cr.assign_memory[463]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[464]= 1'b0;
s.tt.cr.assign_memory[464]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[465]= 1'b1;
s.tt.cr.assign_memory[465]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[466]= 1'b1;
s.tt.cr.assign_memory[466]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[467]= 1'b0;
s.tt.cr.assign_memory[467]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[468]= 1'b0;
s.tt.cr.assign_memory[468]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[469]= 1'b1;
s.tt.cr.assign_memory[469]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[470]= 1'b0;
s.tt.cr.assign_memory[470]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[471]= 1'b1;
s.tt.cr.assign_memory[471]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[472]= 1'b0;
s.tt.cr.assign_memory[472]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[473]= 1'b0;
s.tt.cr.assign_memory[473]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[474]= 1'b1;
s.tt.cr.assign_memory[474]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[475]= 1'b0;
s.tt.cr.assign_memory[475]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[476]= 1'b0;
s.tt.cr.assign_memory[476]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[477]= 1'b0;
s.tt.cr.assign_memory[477]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[478]= 1'b1;
s.tt.cr.assign_memory[478]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[479]= 1'b0;
s.tt.cr.assign_memory[479]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[480]= 1'b1;
s.tt.cr.assign_memory[480]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[481]= 1'b1;
s.tt.cr.assign_memory[481]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[482]= 1'b1;
s.tt.cr.assign_memory[482]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[483]= 1'b1;
s.tt.cr.assign_memory[483]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[484]= 1'b0;
s.tt.cr.assign_memory[484]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[485]= 1'b1;
s.tt.cr.assign_memory[485]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[486]= 1'b1;
s.tt.cr.assign_memory[486]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[487]= 1'b1;
s.tt.cr.assign_memory[487]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[488]= 1'b0;
s.tt.cr.assign_memory[488]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[489]= 1'b1;
s.tt.cr.assign_memory[489]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[490]= 1'b1;
s.tt.cr.assign_memory[490]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[491]= 1'b1;
s.tt.cr.assign_memory[491]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[492]= 1'b1;
s.tt.cr.assign_memory[492]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[493]= 1'b0;
s.tt.cr.assign_memory[493]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[494]= 1'b0;
s.tt.cr.assign_memory[494]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[495]= 1'b0;
s.tt.cr.assign_memory[495]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[496]= 1'b0;
s.tt.cr.assign_memory[496]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[497]= 1'b0;
s.tt.cr.assign_memory[497]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[498]= 1'b1;
s.tt.cr.assign_memory[498]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[499]= 1'b0;
s.tt.cr.assign_memory[499]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[500]= 1'b0;
s.tt.cr.assign_memory[500]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[501]= 1'b0;
s.tt.cr.assign_memory[501]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[502]= 1'b1;
s.tt.cr.assign_memory[502]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[503]= 1'b0;
s.tt.cr.assign_memory[503]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[504]= 1'b0;
s.tt.cr.assign_memory[504]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[505]= 1'b0;
s.tt.cr.assign_memory[505]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[506]= 1'b0;
s.tt.cr.assign_memory[506]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[507]= 1'b0;
s.tt.cr.assign_memory[507]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[508]= 1'b0;
s.tt.cr.assign_memory[508]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[509]= 1'b0;
s.tt.cr.assign_memory[509]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[510]= 1'b0;
s.tt.cr.assign_memory[510]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[511]= 1'b0;
s.tt.cr.assign_memory[511]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[512]= 1'b0;
s.tt.cr.assign_memory[512]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[513]= 1'b0;
s.tt.cr.assign_memory[513]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[514]= 1'b0;
s.tt.cr.assign_memory[514]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[515]= 1'b0;
s.tt.cr.assign_memory[515]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[516]= 1'b0;
s.tt.cr.assign_memory[516]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[517]= 1'b0;
s.tt.cr.assign_memory[517]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[518]= 1'b1;
s.tt.cr.assign_memory[518]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[519]= 1'b0;
s.tt.cr.assign_memory[519]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[520]= 1'b1;
s.tt.cr.assign_memory[520]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[521]= 1'b0;
s.tt.cr.assign_memory[521]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[522]= 1'b0;
s.tt.cr.assign_memory[522]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[523]= 1'b1;
s.tt.cr.assign_memory[523]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[524]= 1'b1;
s.tt.cr.assign_memory[524]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[525]= 1'b0;
s.tt.cr.assign_memory[525]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[526]= 1'b0;
s.tt.cr.assign_memory[526]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[527]= 1'b0;
s.tt.cr.assign_memory[527]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[528]= 1'b1;
s.tt.cr.assign_memory[528]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[529]= 1'b0;
s.tt.cr.assign_memory[529]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[530]= 1'b0;
s.tt.cr.assign_memory[530]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[531]= 1'b1;
s.tt.cr.assign_memory[531]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[532]= 1'b1;
s.tt.cr.assign_memory[532]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[533]= 1'b1;
s.tt.cr.assign_memory[533]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[534]= 1'b1;
s.tt.cr.assign_memory[534]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[535]= 1'b0;
s.tt.cr.assign_memory[535]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[536]= 1'b0;
s.tt.cr.assign_memory[536]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[537]= 1'b0;
s.tt.cr.assign_memory[537]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[538]= 1'b1;
s.tt.cr.assign_memory[538]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[539]= 1'b0;
s.tt.cr.assign_memory[539]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[540]= 1'b1;
s.tt.cr.assign_memory[540]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[541]= 1'b0;
s.tt.cr.assign_memory[541]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[542]= 1'b1;
s.tt.cr.assign_memory[542]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[543]= 1'b1;
s.tt.cr.assign_memory[543]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[544]= 1'b0;
s.tt.cr.assign_memory[544]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[545]= 1'b1;
s.tt.cr.assign_memory[545]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[546]= 1'b0;
s.tt.cr.assign_memory[546]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[547]= 1'b1;
s.tt.cr.assign_memory[547]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[548]= 1'b1;
s.tt.cr.assign_memory[548]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[549]= 1'b1;
s.tt.cr.assign_memory[549]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[550]= 1'b1;
s.tt.cr.assign_memory[550]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[551]= 1'b0;
s.tt.cr.assign_memory[551]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[552]= 1'b1;
s.tt.cr.assign_memory[552]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[553]= 1'b0;
s.tt.cr.assign_memory[553]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[554]= 1'b0;
s.tt.cr.assign_memory[554]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[555]= 1'b1;
s.tt.cr.assign_memory[555]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[556]= 1'b1;
s.tt.cr.assign_memory[556]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[557]= 1'b1;
s.tt.cr.assign_memory[557]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[558]= 1'b0;
s.tt.cr.assign_memory[558]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[559]= 1'b0;
s.tt.cr.assign_memory[559]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[560]= 1'b1;
s.tt.cr.assign_memory[560]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[561]= 1'b0;
s.tt.cr.assign_memory[561]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[562]= 1'b1;
s.tt.cr.assign_memory[562]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[563]= 1'b0;
s.tt.cr.assign_memory[563]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[564]= 1'b1;
s.tt.cr.assign_memory[564]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[565]= 1'b0;
s.tt.cr.assign_memory[565]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[566]= 1'b0;
s.tt.cr.assign_memory[566]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[567]= 1'b1;
s.tt.cr.assign_memory[567]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[568]= 1'b0;
s.tt.cr.assign_memory[568]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[569]= 1'b1;
s.tt.cr.assign_memory[569]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[570]= 1'b0;
s.tt.cr.assign_memory[570]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[571]= 1'b0;
s.tt.cr.assign_memory[571]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[572]= 1'b0;
s.tt.cr.assign_memory[572]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[573]= 1'b1;
s.tt.cr.assign_memory[573]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[574]= 1'b1;
s.tt.cr.assign_memory[574]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[575]= 1'b1;
s.tt.cr.assign_memory[575]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[576]= 1'b1;
s.tt.cr.assign_memory[576]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[577]= 1'b0;
s.tt.cr.assign_memory[577]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[578]= 1'b1;
s.tt.cr.assign_memory[578]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[579]= 1'b0;
s.tt.cr.assign_memory[579]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[580]= 1'b0;
s.tt.cr.assign_memory[580]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[581]= 1'b1;
s.tt.cr.assign_memory[581]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[582]= 1'b1;
s.tt.cr.assign_memory[582]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[583]= 1'b0;
s.tt.cr.assign_memory[583]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[584]= 1'b0;
s.tt.cr.assign_memory[584]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[585]= 1'b0;
s.tt.cr.assign_memory[585]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[586]= 1'b1;
s.tt.cr.assign_memory[586]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[587]= 1'b1;
s.tt.cr.assign_memory[587]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[588]= 1'b0;
s.tt.cr.assign_memory[588]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[589]= 1'b1;
s.tt.cr.assign_memory[589]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[590]= 1'b1;
s.tt.cr.assign_memory[590]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[591]= 1'b0;
s.tt.cr.assign_memory[591]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[592]= 1'b1;
s.tt.cr.assign_memory[592]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[593]= 1'b0;
s.tt.cr.assign_memory[593]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[594]= 1'b0;
s.tt.cr.assign_memory[594]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[595]= 1'b0;
s.tt.cr.assign_memory[595]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[596]= 1'b1;
s.tt.cr.assign_memory[596]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[597]= 1'b0;
s.tt.cr.assign_memory[597]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[598]= 1'b0;
s.tt.cr.assign_memory[598]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[599]= 1'b1;
s.tt.cr.assign_memory[599]= 1'b1;
#`dp_delay_time
s.tt.cr.share_memory[600]= 1'b0;
s.tt.cr.assign_memory[600]= 1'b1;
  
  end
  
  
  
  task print_result;
    for(int i=0;i<`var_num+1;++i) begin
	  $fwrite(fout,"%b\n",s.pe.evaluator2.var_table[i]);
	end
	$fclose(fout);
	
	//$fclose(funsat);
	$display("flip times: %d",s.tt.cr.flip_time);
  
  endtask
  
  
  
endmodule
