`include "clause_evaluator.sv"
module clause_evaluator_array(
  input clk,
  input rst,
  
);

  
  

endmodule